/*
Build a circuit with no inputs and one output. That output should always drive 1 (or logic high).
*/

module top_module( output one );

    // width is 1 bit
    // format is binary
    // value is 1
    assign one = 1'b1

endmodule